-- ######################################################################################################################################################################################################
-- file :
--     gen_heartbeat_wrapper_zedboard.vhd
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     gen_heartbeat.vhd simulation wrapper for ZedBoard evaluation board manufactured by Digilent.
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     register tranfer level (RTL)
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2023-11-11
--         file creation
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01.00. libraries
--     02.00. entity
--     03.00. architecture
--         03.01. components declaration
--             03.01.01. ip_pll
--             03.01.02. gen_heartbeat
--         03.02. signals
--             03.02.01. ip_pll
--             03.02.02. gen_heartbeat
--         03.03. input assignment
--         03.04. components instanciation
--             03.04.01. ip_pll
--             03.04.02. gen_heartbeat
--         03.05. output assignment
-- ######################################################################################################################################################################################################

-- ######################################################################################################################################################################################################
-- 01. libraries
-- ######################################################################################################################################################################################################
    -- ==================================================================================================================================================================================================
	-- 03.01. standard
    -- ==================================================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	
	-- ==================================================================================================================================================================================================
	-- 03.01. custom
    -- ==================================================================================================================================================================================================
    library work;
        use work.pkg_gen_heartbeat_wrapper_zedboard.all;
	
-- ######################################################################################################################################################################################################
-- 02. entity
-- ######################################################################################################################################################################################################

entity gen_heartbeat_wrapper_zedboard is
    port (
	     OSC_100M    : in  std_logic
		;BTNC        : in  std_logic
		;ALIVE       : out std_logic
		;MMCM_LOCKED : out std_logic
		;FAILURE     : out std_logic
	);
end entity gen_heartbeat_wrapper_zedboard;

-- ######################################################################################################################################################################################################
-- 03. architecture
-- ######################################################################################################################################################################################################

architecture schematic of gen_heartbeat_wrapper_zedboard is

    -- ==================================================================================================================================================================================================
	-- 03.01. components declaration
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.01. ip_mmcm
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        component ip_mmcm is
            port (
	             clk_in1  : in  std_logic
		        ;reset    : in  std_logic
				;locked   : out std_logic
				;clk_out1 : out std_logic
	        );
        end component ip_mmcm;
		
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.02. gen_heartbeat
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        component gen_heartbeat is
            generic (
	             g_clk_i_freq : integer
		        ;g_clk_o_freq : integer
	        );
            port (
	             i_clk   : in  std_logic
		        ;i_rst   : in  std_logic
		        ;o_alive : out std_logic
				;o_error : out std_logic_vector(7 downto 0)
	        );
        end component gen_heartbeat;

    -- ==================================================================================================================================================================================================
	-- 03.02. signals
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.01. ip_mmcm
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    signal s_ip_mmcm_i_clk    : std_logic;
	    signal s_ip_mmcm_o_clk    : std_logic;
		signal s_ip_mmcm_i_rst    : std_logic;
	    signal s_ip_mmcm_o_locked : std_logic;
		
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.02. gen_heartbeat
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    signal s_dut_i_rst   : std_logic;
	    signal s_dut_o_alive : std_logic;
		signal s_dut_o_error : std_logic_vector(7 downto 0);
		signal s_error       : std_logic;

begin

    -- ==================================================================================================================================================================================================
	-- 03.03. input assignment
    -- ==================================================================================================================================================================================================
	s_ip_mmcm_i_clk <= OSC_100M;
	s_ip_mmcm_i_rst <= BTNC;

    -- ==================================================================================================================================================================================================
	-- 03.05. DUT reset management
    -- ==================================================================================================================================================================================================
    p_dut_rst_gen : process(s_ip_mmcm_o_locked)
	begin
	    if (s_ip_mmcm_o_locked = '0') then
		    s_dut_i_rst <= '1';
		else
		    s_dut_i_rst <= '0';    
		end if;
	end process p_dut_rst_gen;

    -- ==================================================================================================================================================================================================
	-- 03.05. components instanciation
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.01. ip_mmcm
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_ip_mmcm : ip_mmcm
            port map (
	             clk_in1  => s_ip_mmcm_i_clk
		        ,reset    => s_ip_mmcm_i_rst
				,locked   => s_ip_mmcm_o_locked
				,clk_out1 => s_ip_mmcm_o_clk
	        );

	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.02. DUT : gen_heartbeat
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_dut_gen_heartbeat : gen_heartbeat
            generic map (
	             g_clk_i_freq => c_mmcm_freq
		        ,g_clk_o_freq => c_heartbeat_freq
	        )
            port map (
	             i_clk   => s_ip_mmcm_o_clk
		        ,i_rst   => s_dut_i_rst
		        ,o_alive => s_dut_o_alive
				,o_error => s_dut_o_error
	        );

    -- ==================================================================================================================================================================================================
	-- 03.04. parsing DUT error vector
    -- ==================================================================================================================================================================================================
	p_check_dut_error : process(s_dut_i_rst,s_ip_mmcm_o_clk)
	    variable v_error : std_logic;
	begin
	    if (s_dut_i_rst = '1') then
	        v_error := '0';
			s_error <= '0';
	    elsif (rising_edge(s_ip_mmcm_o_clk)) then
		    v_error := '0';
			-- parsing s_dut_o_error error vector
		    for i in 0 to s_dut_o_error'length-1 loop
		        -- error detected
			    if (s_dut_o_error(i) = '1') then
				    v_error := '1';
				end if;
			end loop;
			s_error <= v_error;
		end if;
	end process p_check_dut_error;	

    -- ==================================================================================================================================================================================================
	-- 03.06. output assignment
    -- ==================================================================================================================================================================================================
	ALIVE       <= s_dut_o_alive;
	MMCM_LOCKED <= s_ip_mmcm_o_locked;
	FAILURE     <= s_error;

end architecture schematic;

-- ######################################################################################################################################################################################################
-- EOF
-- ######################################################################################################################################################################################################