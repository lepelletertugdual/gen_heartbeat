-- ######################################################################################################################################################################################################
-- file :
--     bch_gen_heartbeat_wrapper_zedboard.vhd
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     gen_heartbeat_wrapper_zedboard_sim.vhd testbench file.
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     behavioral
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2022-04-22
--         file creation
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01. libraries
--         01.01. standard
--         01.02. custom
--     02. entity
--     03. architecture
--         03.01. component declaration
--             03.01.01. DUT : gen_heartbeat_wrapper_zedboard_sim
--         03.02. files
--             03.02.01. LOG
--             03.02.02. RPT
--         03.03. constants
--             03.03.01. SIM
--             03.03.02. DUT : gen_heartbeat_wrapper_zedboard_sim
--             03.03.04. files
--         03.04. types
--             03.04.01. FSM
--                 03.04.01.01. fsm_main
--                 03.04.01.02. fsm_init
--                 03.04.01.03. fsm_test
--                 03.04.01.04. fsm_file_mgt_log
--                 03.04.01.05. fsm_file_mgt_rpt
--             03.04.02. test status
--         03.05. signals
--             03.05.01. SIM
--                 03.05.01.01. FSM
--                 03.05.01.02. files
--                 03.05.01.03. clock
--                 03.05.01.04. reset
--                 03.05.01.05. testbench
--             03.05.03. DUT : gen_heartbeat_wrapper_zedboard_sim
--                 03.05.03.01. clock
--                 03.05.03.02. reset
--                 03.05.03.03. indicators
--         03.06. component instanciation
--             03.06.01. DUT : gen_heartbeat_wrapper_zedboard_sim
--         03.07. reinit
--             03.07.01. SIM
--             03.07.02. DUT    
--         03.08. clock generation
--             03.08.01. DUT
--             03.08.02. SIM
--         03.09. fsm_main
--         03.10. fsm_init
--         03.11. fsm_test
--         03.12. fsm_file_mgt_log
--         03.13. fsm_file_mgt_rpt
--         03.14. DUT failure indicator
--         03.15. simulation abort
-- ######################################################################################################################################################################################################

-- ######################################################################################################################################################################################################
-- 01. libraries
-- ######################################################################################################################################################################################################
    -- ==================================================================================================================================================================================================
	-- 01.01. standard
    -- ==================================================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	    use ieee.numeric_std.all;
	    use ieee.math_real.all;
	
    library std;
        use std.textio.all;

    -- ==================================================================================================================================================================================================
	-- 01.02. custom
    -- ==================================================================================================================================================================================================
    library work;
        use work.pkg_mgt_file.all;
		use work.pkg_gen_heartbeat_wrapper_zedboard_sim.all;
	
-- ######################################################################################################################################################################################################
-- 02. entity
-- ######################################################################################################################################################################################################

entity bch_gen_heartbeat_wrapper_zedboard is
end entity bch_gen_heartbeat_wrapper_zedboard;

-- ######################################################################################################################################################################################################
-- 03. architecture
-- ######################################################################################################################################################################################################

architecture behavioral of bch_gen_heartbeat_wrapper_zedboard is

    -- ==================================================================================================================================================================================================
	-- 03.01. component declaration
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.01. DUT : gen_heartbeat_wrapper_zedboard_sim
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        component gen_heartbeat_wrapper_zedboard_sim is
            port (
	            OSC_100M    : in  std_logic
			   ;BTNC        : in  std_logic
		       ;ALIVE       : out std_logic
		       ;MMCM_LOCKED : out std_logic
		       ;FAILURE     : out std_logic
	        );
        end component gen_heartbeat_wrapper_zedboard_sim;

    -- ==================================================================================================================================================================================================
	-- 03.02. files
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.01. LOG
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        file f_file_log : text;

	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.02. RPT
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        file f_file_rpt : text;

    -- ==================================================================================================================================================================================================
	-- 03.03. constants
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. SIM
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_sim_clk_frequency   : integer := 1_000_000_000;
	    constant c_sim_clk_delay       : time    := 0.9 us;
	    constant c_sim_rst_delay       : time    := 0.3 us;
        constant c_sim_clk_period_ns   : time    := integer((real(1)/real(c_sim_clk_frequency))*1.0e9)*1 ns;
	    constant c_sim_clk_period      : real    := real(1)/real(c_sim_clk_frequency);
	
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.02. DUT : gen_heartbeat_wrapper_zedboard_sim
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_osc_delay        : time    := 2.4 us;
	    constant c_dut_rst_delay    : time    := 1.3 us;
        constant c_osc_period_ns    : time    := integer((real(1)/real(c_osc_freq))*1.0e9)*1 ns;
	    constant c_dut_clk_period   : real    := real(1)/real(c_osc_freq);
	    constant c_heartbeat_period : real    := real(1)/real(c_heartbeat_freq);
	    constant c_alive_cycle_full : integer := integer(real(c_heartbeat_period)/real(c_sim_clk_period));
	    constant c_alive_cycle_half : integer := integer(real(c_alive_cycle_full)/real(2));
	
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.03. simulation duration
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		constant c_sim_duration_factor : integer := 16;
	    constant c_sim_duration_ns     : integer := integer(real(c_sim_duration_factor)*real(c_heartbeat_period)/real(c_sim_clk_period));
	
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.03. file
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		constant c_file_log_name : string := "log_bch_gen_heartbeat_wrapper_zedboard.csv";
		constant c_file_rpt_name : string := "rpt_bch_gen_heartbeat_wrapper_zedboard.txt";
	
    -- ==================================================================================================================================================================================================
	-- 03.04. types
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.01. FSM
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- ==========================================================================================================================================================================================
			-- 03.04.01.01. fsm_main
			-- ==========================================================================================================================================================================================
	        type t_fsm_main is (
	             state_fsm_main_start
                ,state_fsm_main_file_rpt_open
                ,state_fsm_main_file_log_open
			    ,state_fsm_main_init
		        ,state_fsm_main_run
                ,state_fsm_main_file_rpt_close
                ,state_fsm_main_file_log_close
		        ,state_fsm_main_stop
	        );

		    -- ==========================================================================================================================================================================================
			-- 03.04.01.02. fsm_init
			-- ==========================================================================================================================================================================================
	        type t_fsm_init is (
	             state_fsm_init_idle
		        ,state_fsm_init_run
		        ,state_fsm_init_done
	        );

		    -- ==========================================================================================================================================================================================
			-- 03.04.01.03. fsm_test
			-- ==========================================================================================================================================================================================
	        type t_fsm_test is (
	             state_fsm_test_idle
		        ,state_fsm_test_run
		        ,state_fsm_test_done
	        );
	
		    -- ==========================================================================================================================================================================================
			-- 03.04.01.04. fsm_file_mgt_log
			-- ==========================================================================================================================================================================================
	        type t_fsm_file_mgt_log is (
	             state_fsm_file_mgt_log_open
				,state_fsm_file_mgt_log_write_head
	            ,state_fsm_file_mgt_log_write_data
		        ,state_fsm_file_mgt_log_close
				,state_fsm_file_mgt_log_done
	        );

		    -- ==========================================================================================================================================================================================
			-- 03.04.01.04. fsm_file_mgt_rpt
			-- ==========================================================================================================================================================================================
	        type t_fsm_file_mgt_rpt is (
	             state_fsm_file_mgt_rpt_open
	            ,state_fsm_file_mgt_rpt_write_status
		        ,state_fsm_file_mgt_rpt_close
				,state_fsm_file_mgt_rpt_done
	        );

	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.02. test status
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	        type t_sim_test_status is (
	             TEST_OK
	            ,TEST_KO
	        );
	
    -- ==================================================================================================================================================================================================
	-- 03.05. signals
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.02. SIM
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- ==========================================================================================================================================================================================
			-- 03.05.02.01. FSM
			-- ==========================================================================================================================================================================================
	        signal s_fsm_main_state   : t_fsm_main;
	        signal s_fsm_init_state   : t_fsm_init;
	        signal s_fsm_test_state   : t_fsm_test;
		    signal s_fsm_file_mgt_log : t_fsm_file_mgt_log;
		    signal s_fsm_file_mgt_rpt : t_fsm_file_mgt_rpt;
	
		    -- ==========================================================================================================================================================================================
			-- 03.05.02.02. files
			-- ==========================================================================================================================================================================================
		    signal s_sim_file_req_log_open  : std_logic;
		    signal s_sim_file_ack_log_open  : std_logic;
		    signal s_sim_file_req_log_close : std_logic;
		    signal s_sim_file_ack_log_close : std_logic;
		    signal s_sim_file_req_rpt_open  : std_logic;
		    signal s_sim_file_ack_rpt_open  : std_logic;
		    signal s_sim_file_req_rpt_close : std_logic;
		    signal s_sim_file_ack_rpt_close : std_logic;
			
		    -- ==========================================================================================================================================================================================
			-- 03.05.02.03. clock
			-- ==========================================================================================================================================================================================
            signal s_sim_clk : std_logic;
			
		    -- ==========================================================================================================================================================================================
			-- 03.05.02.04. reset
			-- ==========================================================================================================================================================================================
		    signal s_sim_rst : std_logic;
			
		    -- ==========================================================================================================================================================================================
			-- 03.05.02.05. testbench
			-- ==========================================================================================================================================================================================
	        signal s_sim_cnt         : integer range 0 to c_sim_duration_ns-1;
		    signal s_sim_done        : std_logic;
		    signal s_sim_init_req    : std_logic;
		    signal s_sim_init_ack    : std_logic;
		    signal s_sim_test_req    : std_logic;
		    signal s_sim_test_ack    : std_logic;
		    signal s_sim_test_status : t_sim_test_status;
	
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.03. DUT : gen_heartbeat_wrapper_zedboard_sim
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- ==========================================================================================================================================================================================
			-- 03.05.03.01. clock
			-- ==========================================================================================================================================================================================
	        signal s_dut_i_osc : std_logic;
			
		    -- ==========================================================================================================================================================================================
			-- 03.05.03.02. reset
			-- ==========================================================================================================================================================================================
	        signal s_dut_i_rst : std_logic;
			
		    -- ==========================================================================================================================================================================================
			-- 03.05.03.03. indicators
			-- ==========================================================================================================================================================================================			
		    signal s_dut_o_alive       : std_logic;
		    signal s_dut_o_mmcm_locked : std_logic;
		    signal s_dut_o_failure     : std_logic;

begin

    -- ==================================================================================================================================================================================================
	-- 03.06. component instanciation
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.01. DUT : gen_heartbeat_wrapper_zedboard_sim
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_dut_gen_heartbeat_wrapper_zedboard_sim : gen_heartbeat_wrapper_zedboard_sim
            port map (
	             OSC_100M    => s_dut_i_osc
				,BTNC        => s_dut_i_rst
		        ,ALIVE       => s_dut_o_alive
		        ,MMCM_LOCKED => s_dut_o_mmcm_locked
		        ,FAILURE     => s_dut_o_failure
	        );

    -- ==================================================================================================================================================================================================
	-- 03.07. reinit
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.01. SIM reinit
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_sim_rst   <= '1','0' after c_sim_rst_delay;

	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.01. DUT reinit
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_dut_i_rst <= '1','0' after c_dut_rst_delay;

    -- ==================================================================================================================================================================================================
	-- 03.08. clock generation
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.08.01. SIM
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_sim_clk : process
		begin
	        s_sim_clk <= '0';
	        wait for c_sim_clk_delay;
		    while true loop
		        s_sim_clk <= '1';
			    wait for c_sim_clk_period_ns/2;
			    s_sim_clk <= '0';
			    wait for c_sim_clk_period_ns/2;
		    end loop;
	    end process p_gen_sim_clk;

	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.08.02. DUT
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_osc : process
		begin
	        s_dut_i_osc <= '0';
	        wait for c_osc_delay;
		    while true loop
		        s_dut_i_osc <= '1';
			    wait for c_osc_period_ns/2;
			    s_dut_i_osc <= '0';
			    wait for c_osc_period_ns/2;
		    end loop;
	    end process p_gen_osc;

    -- ==================================================================================================================================================================================================
	-- 03.09. fsm_main
    -- ==================================================================================================================================================================================================
	p_fsm_main : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_main_state <= state_fsm_main_start;
			s_sim_done <= '0';
			s_sim_init_req <= '0';
			s_sim_test_req <= '0';
			s_sim_file_req_log_open <= '0';
			s_sim_file_req_log_close <= '0';
			s_sim_file_req_rpt_open <= '0';
			s_sim_file_req_rpt_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_done <= '0';
            s_sim_init_req <= '0';
			s_sim_test_req <= '0';
			s_sim_file_req_log_open <= '0';
			s_sim_file_req_log_close <= '0';
			s_sim_file_req_rpt_open <= '0';
			s_sim_file_req_rpt_close <= '0';
		    case s_fsm_main_state is
			    -- wait for DUT clock locking
				when state_fsm_main_start =>
				    if (s_dut_o_mmcm_locked = '1') then
					    s_fsm_main_state <= state_fsm_main_file_rpt_open;
						s_sim_file_req_rpt_open <= '1';
					end if;
				-- wait for RPT file to be opened
			    when state_fsm_main_file_rpt_open =>
				    if (s_sim_file_ack_rpt_open = '1') then
					    s_fsm_main_state <= state_fsm_main_file_log_open;
					    s_sim_file_req_log_open <= '1';
					end if;
				-- wait for LOG file to be opened
				when state_fsm_main_file_log_open =>
				    if (s_sim_file_ack_log_open = '1') then
					    s_fsm_main_state <= state_fsm_main_init;
						s_sim_init_req <= '1';
					end if;
				-- waiting for init done
				when state_fsm_main_init =>
				    if (s_sim_init_ack = '1') then
					    s_fsm_main_state <= state_fsm_main_run;
					    s_sim_test_req <= '1';
					end if;
				-- waiting for test done
				when state_fsm_main_run =>
                    if (s_sim_test_ack = '1') then
					    s_fsm_main_state <= state_fsm_main_file_log_close;
						s_sim_file_req_log_close <= '1';
					end if;
				-- waiting for data file to be closed
				when state_fsm_main_file_log_close =>
                    if (s_sim_file_ack_log_close = '1') then
					    s_fsm_main_state <= state_fsm_main_file_rpt_close;
						s_sim_file_req_rpt_close <= '1';
					end if;
				-- waiting for SIM report file to be closed
				when state_fsm_main_file_rpt_close =>
                    if (s_sim_file_ack_rpt_close = '1') then
					    s_fsm_main_state <= state_fsm_main_stop;
				        s_sim_done <= '1';
					end if;
				-- test stopped
                when state_fsm_main_stop =>
                    null;
			end case;
		end if;
	end process p_fsm_main;

    -- ==================================================================================================================================================================================================
	-- 03.10. fsm_init
    -- ==================================================================================================================================================================================================
	fsm_init : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_init_state <= state_fsm_init_idle;
			s_sim_init_ack <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_init_ack <= '0';
		    case s_fsm_init_state is
			    -- waiting for init request
			    when state_fsm_init_idle =>
				    if (s_sim_init_req = '1') then
					    s_fsm_init_state <= state_fsm_init_run;
					end if;
				-- running init
				when state_fsm_init_run =>
					s_fsm_init_state <= state_fsm_init_done;
                    s_sim_init_ack <= '1';
				-- init done
                when state_fsm_init_done =>
				    null;
			end case;
		end if;
	end process fsm_init;

    -- ==================================================================================================================================================================================================
	-- 03.11. fsm_test
    -- ==================================================================================================================================================================================================
	p_fsm_test : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_test_state <= state_fsm_test_idle;
			s_sim_cnt <= 0;
			s_sim_test_ack <= '0';
			s_sim_test_status <= TEST_OK;
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_test_ack <= '0';
		    case s_fsm_test_state is
			    -- waiting for test request
			    when state_fsm_test_idle =>
				    if (s_sim_test_req = '1') then
					    s_fsm_test_state <= state_fsm_test_run;
					end if;
				-- running test
				when state_fsm_test_run =>
				    if (s_sim_cnt = c_sim_duration_ns-1) then
					    s_sim_test_ack <= '1';
					    s_fsm_test_state <= state_fsm_test_done;
					    s_sim_cnt <= 0;
						s_sim_test_status <= TEST_OK;
                    else
					    s_sim_cnt <= s_sim_cnt + 1;
					end if;
				-- test done
                when state_fsm_test_done =>
                    null;
			end case;
		end if;
	end process p_fsm_test;

    -- ==================================================================================================================================================================================================
	-- 03.12. fsm_file_mgt_log
    -- ==================================================================================================================================================================================================
	p_fsm_file_mgt_log : process(s_sim_rst,s_sim_clk)
		constant c_justified  : side   := right;
		constant c_field      : width  := 0;
		constant c_unit       : time   := ns;
		constant c_separator  : string := ",";
		constant c_value_head : string := "time,data";
	    variable v_value_time : time;
		variable v_value_data : string(1 to 4);
		variable v_value_foot : string(1 to 7);
		variable v_line       : line;
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_open;
		    s_sim_file_ack_log_open <= '0';
			s_sim_file_ack_log_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_file_ack_log_open <= '0';
			s_sim_file_ack_log_close <= '0';
            case s_fsm_file_mgt_log is
                -- open file
			    when state_fsm_file_mgt_log_open =>
				    if (s_sim_file_req_log_open = '1') then
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_write_head;
						s_sim_file_ack_log_open <= '1';
						proc_file_log_open(c_file_log_name,f_file_log);
					end if;
				-- write header
				when state_fsm_file_mgt_log_write_head =>
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_write_data;
						write(v_line,c_value_head,c_justified,c_field);
	                    writeline(f_file_log,v_line);
				-- write data
				when state_fsm_file_mgt_log_write_data =>
				    if (s_sim_file_req_log_close = '1') then
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_close;
						-- timestamp
						v_value_time := now;
						write(v_line,v_value_time,c_justified,c_field,c_unit);
						-- separator
						write(v_line,c_separator,c_justified,c_field);
						-- data value
						v_value_data := "NONE";
					    write(v_line,v_value_data,c_justified,c_field);
	                    writeline(f_file_log,v_line);
					end if;
                -- close file
				when state_fsm_file_mgt_log_close =>
					s_fsm_file_mgt_log <= state_fsm_file_mgt_log_done;
				    s_sim_file_ack_log_close <= '1';
                    proc_file_log_close(c_file_log_name,f_file_log);
				-- done
				when state_fsm_file_mgt_log_done  =>
				    null;
			end case;
		end if;
	end process p_fsm_file_mgt_log;

    -- ==================================================================================================================================================================================================
	-- 03.13. fsm_file_mgt_rpt
    -- ==================================================================================================================================================================================================
	p_fsm_file_mgt_rpt : process(s_sim_rst,s_sim_clk)
		constant c_justified    : side  := right;
		constant c_field        : width := 0;
		variable v_value_status : string(1 to 7);
		variable v_line         : line;
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_open;
		    s_sim_file_ack_rpt_open <= '0';
			s_sim_file_ack_rpt_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_file_ack_rpt_open <= '0';
			s_sim_file_ack_rpt_close <= '0';
            case s_fsm_file_mgt_rpt is
                -- open file
			    when state_fsm_file_mgt_rpt_open =>
				    if (s_sim_file_req_rpt_open = '1') then
					    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_write_status;
						s_sim_file_ack_rpt_open <= '1';
						proc_file_rpt_open(c_file_rpt_name,f_file_rpt);
					end if;
				-- write status
				when state_fsm_file_mgt_rpt_write_status =>
				    if (s_sim_file_req_rpt_close = '1') then
					    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_close;
					    -- write test status
					    case s_sim_test_status is
					        when TEST_OK => v_value_status := "TEST_OK";
						    when others  => v_value_status := "TEST_KO";
					    end case;
					    write(v_line,v_value_status,c_justified,c_field);
	                    writeline(f_file_rpt,v_line);
					end if;
                -- close file
				when state_fsm_file_mgt_rpt_close =>
					s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_done;
				    s_sim_file_ack_rpt_close <= '1';
                    proc_file_rpt_close(c_file_rpt_name,f_file_rpt);
				-- done
				when state_fsm_file_mgt_rpt_done  =>
				    null;
			end case;
		end if;
	end process p_fsm_file_mgt_rpt;

    -- ==================================================================================================================================================================================================
	-- 03.14. DUT failure indicator
    -- ==================================================================================================================================================================================================
	p_sim_abort_default : process(s_sim_clk)
	begin
	    if (rising_edge(s_sim_clk)) then
		    if (s_dut_o_failure = '1') then
		        assert false
			        report "end of simulation - DUT failure : default detected" 
		 	            severity failure;
			end if;
		end if;
	end process p_sim_abort_default;

    -- ==================================================================================================================================================================================================
	-- 03.15. simulation abort
    -- ==================================================================================================================================================================================================
	p_sim_abort_nominal : process(s_sim_clk)
	begin
		if (rising_edge(s_sim_clk)) then
            if (s_sim_done = '1') then
			    assert false 
				    report "end of simulation - success" 
					    severity failure;
			end if;
		end if;
	end process p_sim_abort_nominal;

end architecture behavioral;

-- ######################################################################################################################################################################################################
-- EOF
-- ######################################################################################################################################################################################################